module cpu_2601 (
    /* verilator lint_off UNUSED */
    input  logic clk,
    input  logic rst
    /* verilator lint_on UNUSED */
);


endmodule
